library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity mlp_rom is
    Port (
        addr : in integer range 0 to 2345;
        data_out : out signed(8 downto 0) -- Q1.8 format
    );
end mlp_rom;

architecture Behavioral of mlp_rom is
    type rom_array is array (0 to 2345) of signed(8 downto 0); -- 1984 + 320 + 32 + 10
    
    signal rom : rom_array := (

    -- weights_L2 - 1984 addresses (hidden layer weights):
    0 => to_signed(-41, 9),
    1 => to_signed(-2, 9),
    2 => to_signed(-5, 9),
    3 => to_signed(0, 9),
    4 => to_signed(-31, 9),
    5 => to_signed(0, 9),
    6 => to_signed(2, 9),
    7 => to_signed(-18, 9),
    8 => to_signed(-30, 9),
    9 => to_signed(-54, 9),
    10 => to_signed(-57, 9),
    11 => to_signed(20, 9),
    12 => to_signed(-7, 9),
    13 => to_signed(-7, 9),
    14 => to_signed(3, 9),
    15 => to_signed(24, 9),
    16 => to_signed(46, 9),
    17 => to_signed(34, 9),
    18 => to_signed(-12, 9),
    19 => to_signed(0, 9),
    20 => to_signed(-16, 9),
    21 => to_signed(-2, 9),
    22 => to_signed(1, 9),
    23 => to_signed(16, 9),
    24 => to_signed(13, 9),
    25 => to_signed(63, 9),
    26 => to_signed(5, 9),
    27 => to_signed(-25, 9),
    28 => to_signed(-15, 9),
    29 => to_signed(3, 9),
    30 => to_signed(0, 9),
    31 => to_signed(-6, 9),
    32 => to_signed(8, 9),
    33 => to_signed(34, 9),
    34 => to_signed(10, 9),
    35 => to_signed(-28, 9),
    36 => to_signed(-22, 9),
    37 => to_signed(3, 9),
    38 => to_signed(4, 9),
    39 => to_signed(9, 9),
    40 => to_signed(74, 9),
    41 => to_signed(33, 9),
    42 => to_signed(52, 9),
    43 => to_signed(19, 9),
    44 => to_signed(12, 9),
    45 => to_signed(3, 9),
    46 => to_signed(0, 9),
    47 => to_signed(-12, 9),
    48 => to_signed(29, 9),
    49 => to_signed(-22, 9),
    50 => to_signed(14, 9),
    51 => to_signed(27, 9),
    52 => to_signed(8, 9),
    53 => to_signed(3, 9),
    54 => to_signed(-1, 9),
    55 => to_signed(-16, 9),
    56 => to_signed(-28, 9),
    57 => to_signed(7, 9),
    58 => to_signed(14, 9),
    59 => to_signed(4, 9),
    60 => to_signed(-10, 9),
    61 => to_signed(-1, 9),
    62 => to_signed(2, 9),
    63 => to_signed(38, 9),
    64 => to_signed(14, 9),
    65 => to_signed(-25, 9),
    66 => to_signed(-22, 9),
    67 => to_signed(-11, 9),
    68 => to_signed(3, 9),
    69 => to_signed(33, 9),
    70 => to_signed(70, 9),
    71 => to_signed(-13, 9),
    72 => to_signed(7, 9),
    73 => to_signed(17, 9),
    74 => to_signed(-5, 9),
    75 => to_signed(-1, 9),
    76 => to_signed(-1, 9),
    77 => to_signed(1, 9),
    78 => to_signed(-3, 9),
    79 => to_signed(-61, 9),
    80 => to_signed(1, 9),
    81 => to_signed(47, 9),
    82 => to_signed(11, 9),
    83 => to_signed(-2, 9),
    84 => to_signed(3, 9),
    85 => to_signed(-2, 9),
    86 => to_signed(-17, 9),
    87 => to_signed(0, 9),
    88 => to_signed(17, 9),
    89 => to_signed(-21, 9),
    90 => to_signed(-17, 9),
    91 => to_signed(0, 9),
    92 => to_signed(-2, 9),
    93 => to_signed(-6, 9),
    94 => to_signed(-22, 9),
    95 => to_signed(-4, 9),
    96 => to_signed(-7, 9),
    97 => to_signed(-30, 9),
    98 => to_signed(-13, 9),
    99 => to_signed(-1, 9),
    100 => to_signed(-3, 9),
    101 => to_signed(-5, 9),
    102 => to_signed(-9, 9),
    103 => to_signed(-43, 9),
    104 => to_signed(-42, 9),
    105 => to_signed(14, 9),
    106 => to_signed(1, 9),
    107 => to_signed(0, 9),
    108 => to_signed(-3, 9),
    109 => to_signed(9, 9),
    110 => to_signed(40, 9),
    111 => to_signed(10, 9),
    112 => to_signed(-28, 9),
    113 => to_signed(33, 9),
    114 => to_signed(5, 9),
    115 => to_signed(-3, 9),
    116 => to_signed(0, 9),
    117 => to_signed(4, 9),
    118 => to_signed(21, 9),
    119 => to_signed(56, 9),
    120 => to_signed(6, 9),
    121 => to_signed(-9, 9),
    122 => to_signed(-11, 9),
    123 => to_signed(-12, 9),
    124 => to_signed(26, 9),
    125 => to_signed(0, 9),
    126 => to_signed(15, 9),
    127 => to_signed(56, 9),
    128 => to_signed(34, 9),
    129 => to_signed(16, 9),
    130 => to_signed(3, 9),
    131 => to_signed(15, 9),
    132 => to_signed(22, 9),
    133 => to_signed(27, 9),
    134 => to_signed(4, 9),
    135 => to_signed(11, 9),
    136 => to_signed(-2, 9),
    137 => to_signed(6, 9),
    138 => to_signed(0, 9),
    139 => to_signed(11, 9),
    140 => to_signed(19, 9),
    141 => to_signed(-41, 9),
    142 => to_signed(-44, 9),
    143 => to_signed(-35, 9),
    144 => to_signed(-27, 9),
    145 => to_signed(5, 9),
    146 => to_signed(1, 9),
    147 => to_signed(14, 9),
    148 => to_signed(34, 9),
    149 => to_signed(18, 9),
    150 => to_signed(6, 9),
    151 => to_signed(11, 9),
    152 => to_signed(21, 9),
    153 => to_signed(0, 9),
    154 => to_signed(0, 9),
    155 => to_signed(16, 9),
    156 => to_signed(16, 9),
    157 => to_signed(30, 9),
    158 => to_signed(40, 9),
    159 => to_signed(32, 9),
    160 => to_signed(26, 9),
    161 => to_signed(-1, 9),
    162 => to_signed(0, 9),
    163 => to_signed(6, 9),
    164 => to_signed(-34, 9),
    165 => to_signed(7, 9),
    166 => to_signed(15, 9),
    167 => to_signed(0, 9),
    168 => to_signed(-1, 9),
    169 => to_signed(-4, 9),
    170 => to_signed(1, 9),
    171 => to_signed(2, 9),
    172 => to_signed(-38, 9),
    173 => to_signed(-21, 9),
    174 => to_signed(-25, 9),
    175 => to_signed(-44, 9),
    176 => to_signed(-13, 9),
    177 => to_signed(1, 9),
    178 => to_signed(1, 9),
    179 => to_signed(-1, 9),
    180 => to_signed(5, 9),
    181 => to_signed(-9, 9),
    182 => to_signed(-43, 9),
    183 => to_signed(-41, 9),
    184 => to_signed(-20, 9),
    185 => to_signed(-4, 9),
    186 => to_signed(-3, 9),
    187 => to_signed(-1, 9),
    188 => to_signed(-1, 9),
    189 => to_signed(3, 9),
    190 => to_signed(1, 9),
    191 => to_signed(0, 9),
    192 => to_signed(-1, 9),
    193 => to_signed(4, 9),
    194 => to_signed(-4, 9),
    195 => to_signed(2, 9),
    196 => to_signed(0, 9),
    197 => to_signed(-1, 9),
    198 => to_signed(0, 9),
    199 => to_signed(2, 9),
    200 => to_signed(-2, 9),
    201 => to_signed(-5, 9),
    202 => to_signed(0, 9),
    203 => to_signed(-1, 9),
    204 => to_signed(0, 9),
    205 => to_signed(0, 9),
    206 => to_signed(3, 9),
    207 => to_signed(1, 9),
    208 => to_signed(-1, 9),
    209 => to_signed(-1, 9),
    210 => to_signed(-3, 9),
    211 => to_signed(2, 9),
    212 => to_signed(-2, 9),
    213 => to_signed(-4, 9),
    214 => to_signed(-5, 9),
    215 => to_signed(-1, 9),
    216 => to_signed(4, 9),
    217 => to_signed(1, 9),
    218 => to_signed(0, 9),
    219 => to_signed(-2, 9),
    220 => to_signed(-3, 9),
    221 => to_signed(0, 9),
    222 => to_signed(1, 9),
    223 => to_signed(1, 9),
    224 => to_signed(-1, 9),
    225 => to_signed(-2, 9),
    226 => to_signed(0, 9),
    227 => to_signed(0, 9),
    228 => to_signed(-1, 9),
    229 => to_signed(1, 9),
    230 => to_signed(-2, 9),
    231 => to_signed(-1, 9),
    232 => to_signed(1, 9),
    233 => to_signed(2, 9),
    234 => to_signed(-6, 9),
    235 => to_signed(1, 9),
    236 => to_signed(-2, 9),
    237 => to_signed(4, 9),
    238 => to_signed(-3, 9),
    239 => to_signed(3, 9),
    240 => to_signed(-3, 9),
    241 => to_signed(0, 9),
    242 => to_signed(0, 9),
    243 => to_signed(1, 9),
    244 => to_signed(0, 9),
    245 => to_signed(1, 9),
    246 => to_signed(0, 9),
    247 => to_signed(-3, 9),
    248 => to_signed(2, 9),
    249 => to_signed(21, 9),
    250 => to_signed(15, 9),
    251 => to_signed(17, 9),
    252 => to_signed(16, 9),
    253 => to_signed(-7, 9),
    254 => to_signed(0, 9),
    255 => to_signed(15, 9),
    256 => to_signed(28, 9),
    257 => to_signed(20, 9),
    258 => to_signed(32, 9),
    259 => to_signed(23, 9),
    260 => to_signed(-1, 9),
    261 => to_signed(-1, 9),
    262 => to_signed(0, 9),
    263 => to_signed(-3, 9),
    264 => to_signed(-10, 9),
    265 => to_signed(-10, 9),
    266 => to_signed(-3, 9),
    267 => to_signed(19, 9),
    268 => to_signed(17, 9),
    269 => to_signed(1, 9),
    270 => to_signed(-2, 9),
    271 => to_signed(-6, 9),
    272 => to_signed(-7, 9),
    273 => to_signed(-28, 9),
    274 => to_signed(0, 9),
    275 => to_signed(-8, 9),
    276 => to_signed(-32, 9),
    277 => to_signed(4, 9),
    278 => to_signed(2, 9),
    279 => to_signed(-3, 9),
    280 => to_signed(-8, 9),
    281 => to_signed(4, 9),
    282 => to_signed(-17, 9),
    283 => to_signed(-13, 9),
    284 => to_signed(-16, 9),
    285 => to_signed(0, 9),
    286 => to_signed(-6, 9),
    287 => to_signed(-26, 9),
    288 => to_signed(-20, 9),
    289 => to_signed(-36, 9),
    290 => to_signed(-25, 9),
    291 => to_signed(20, 9),
    292 => to_signed(16, 9),
    293 => to_signed(-3, 9),
    294 => to_signed(0, 9),
    295 => to_signed(-22, 9),
    296 => to_signed(10, 9),
    297 => to_signed(-1, 9),
    298 => to_signed(16, 9),
    299 => to_signed(38, 9),
    300 => to_signed(-10, 9),
    301 => to_signed(-7, 9),
    302 => to_signed(2, 9),
    303 => to_signed(5, 9),
    304 => to_signed(14, 9),
    305 => to_signed(56, 9),
    306 => to_signed(27, 9),
    307 => to_signed(-8, 9),
    308 => to_signed(-8, 9),
    309 => to_signed(-5, 9),
    310 => to_signed(22, 9),
    311 => to_signed(19, 9),
    312 => to_signed(30, 9),
    313 => to_signed(41, 9),
    314 => to_signed(17, 9),
    315 => to_signed(2, 9),
    316 => to_signed(-6, 9),
    317 => to_signed(13, 9),
    318 => to_signed(28, 9),
    319 => to_signed(35, 9),
    320 => to_signed(18, 9),
    321 => to_signed(9, 9),
    322 => to_signed(-16, 9),
    323 => to_signed(0, 9),
    324 => to_signed(-1, 9),
    325 => to_signed(-2, 9),
    326 => to_signed(-25, 9),
    327 => to_signed(-19, 9),
    328 => to_signed(-16, 9),
    329 => to_signed(-37, 9),
    330 => to_signed(-22, 9),
    331 => to_signed(-1, 9),
    332 => to_signed(0, 9),
    333 => to_signed(-5, 9),
    334 => to_signed(-16, 9),
    335 => to_signed(2, 9),
    336 => to_signed(20, 9),
    337 => to_signed(-26, 9),
    338 => to_signed(-26, 9),
    339 => to_signed(0, 9),
    340 => to_signed(-1, 9),
    341 => to_signed(-12, 9),
    342 => to_signed(-14, 9),
    343 => to_signed(28, 9),
    344 => to_signed(1, 9),
    345 => to_signed(-13, 9),
    346 => to_signed(-3, 9),
    347 => to_signed(-4, 9),
    348 => to_signed(-3, 9),
    349 => to_signed(-26, 9),
    350 => to_signed(-23, 9),
    351 => to_signed(-13, 9),
    352 => to_signed(-1, 9),
    353 => to_signed(-8, 9),
    354 => to_signed(15, 9),
    355 => to_signed(4, 9),
    356 => to_signed(0, 9),
    357 => to_signed(-9, 9),
    358 => to_signed(7, 9),
    359 => to_signed(3, 9),
    360 => to_signed(18, 9),
    361 => to_signed(18, 9),
    362 => to_signed(-10, 9),
    363 => to_signed(1, 9),
    364 => to_signed(1, 9),
    365 => to_signed(5, 9),
    366 => to_signed(33, 9),
    367 => to_signed(41, 9),
    368 => to_signed(-2, 9),
    369 => to_signed(-19, 9),
    370 => to_signed(-10, 9),
    371 => to_signed(-1, 9),
    372 => to_signed(4, 9),
    373 => to_signed(22, 9),
    374 => to_signed(-9, 9),
    375 => to_signed(-25, 9),
    376 => to_signed(-13, 9),
    377 => to_signed(-6, 9),
    378 => to_signed(-2, 9),
    379 => to_signed(2, 9),
    380 => to_signed(42, 9),
    381 => to_signed(1, 9),
    382 => to_signed(-38, 9),
    383 => to_signed(19, 9),
    384 => to_signed(11, 9),
    385 => to_signed(0, 9),
    386 => to_signed(-3, 9),
    387 => to_signed(-3, 9),
    388 => to_signed(52, 9),
    389 => to_signed(-5, 9),
    390 => to_signed(-34, 9),
    391 => to_signed(90, 9),
    392 => to_signed(30, 9),
    393 => to_signed(0, 9),
    394 => to_signed(-2, 9),
    395 => to_signed(12, 9),
    396 => to_signed(41, 9),
    397 => to_signed(0, 9),
    398 => to_signed(-23, 9),
    399 => to_signed(50, 9),
    400 => to_signed(23, 9),
    401 => to_signed(-2, 9),
    402 => to_signed(-3, 9),
    403 => to_signed(23, 9),
    404 => to_signed(16, 9),
    405 => to_signed(-14, 9),
    406 => to_signed(-30, 9),
    407 => to_signed(-40, 9),
    408 => to_signed(9, 9),
    409 => to_signed(3, 9),
    410 => to_signed(0, 9),
    411 => to_signed(13, 9),
    412 => to_signed(15, 9),
    413 => to_signed(-46, 9),
    414 => to_signed(-25, 9),
    415 => to_signed(0, 9),
    416 => to_signed(1, 9),
    417 => to_signed(0, 9),
    418 => to_signed(-3, 9),
    419 => to_signed(-7, 9),
    420 => to_signed(29, 9),
    421 => to_signed(-5, 9),
    422 => to_signed(-18, 9),
    423 => to_signed(-13, 9),
    424 => to_signed(-12, 9),
    425 => to_signed(-2, 9),
    426 => to_signed(2, 9),
    427 => to_signed(-4, 9),
    428 => to_signed(-5, 9),
    429 => to_signed(46, 9),
    430 => to_signed(22, 9),
    431 => to_signed(-41, 9),
    432 => to_signed(-25, 9),
    433 => to_signed(-12, 9),
    434 => to_signed(13, 9),
    435 => to_signed(37, 9),
    436 => to_signed(-21, 9),
    437 => to_signed(14, 9),
    438 => to_signed(-13, 9),
    439 => to_signed(-8, 9),
    440 => to_signed(-3, 9),
    441 => to_signed(1, 9),
    442 => to_signed(27, 9),
    443 => to_signed(-18, 9),
    444 => to_signed(2, 9),
    445 => to_signed(16, 9),
    446 => to_signed(-18, 9),
    447 => to_signed(-6, 9),
    448 => to_signed(2, 9),
    449 => to_signed(29, 9),
    450 => to_signed(18, 9),
    451 => to_signed(48, 9),
    452 => to_signed(50, 9),
    453 => to_signed(13, 9),
    454 => to_signed(-1, 9),
    455 => to_signed(3, 9),
    456 => to_signed(-2, 9),
    457 => to_signed(-18, 9),
    458 => to_signed(-7, 9),
    459 => to_signed(20, 9),
    460 => to_signed(19, 9),
    461 => to_signed(10, 9),
    462 => to_signed(-46, 9),
    463 => to_signed(2, 9),
    464 => to_signed(3, 9),
    465 => to_signed(-30, 9),
    466 => to_signed(-33, 9),
    467 => to_signed(6, 9),
    468 => to_signed(-11, 9),
    469 => to_signed(-24, 9),
    470 => to_signed(-56, 9),
    471 => to_signed(0, 9),
    472 => to_signed(-2, 9),
    473 => to_signed(-21, 9),
    474 => to_signed(-18, 9),
    475 => to_signed(0, 9),
    476 => to_signed(7, 9),
    477 => to_signed(-34, 9),
    478 => to_signed(-33, 9),
    479 => to_signed(0, 9),
    480 => to_signed(-2, 9),
    481 => to_signed(6, 9),
    482 => to_signed(12, 9),
    483 => to_signed(-14, 9),
    484 => to_signed(20, 9),
    485 => to_signed(-7, 9),
    486 => to_signed(6, 9),
    487 => to_signed(4, 9),
    488 => to_signed(-1, 9),
    489 => to_signed(5, 9),
    490 => to_signed(20, 9),
    491 => to_signed(51, 9),
    492 => to_signed(13, 9),
    493 => to_signed(18, 9),
    494 => to_signed(27, 9),
    495 => to_signed(16, 9),
    496 => to_signed(-6, 9),
    497 => to_signed(20, 9),
    498 => to_signed(24, 9),
    499 => to_signed(18, 9),
    500 => to_signed(-5, 9),
    501 => to_signed(-4, 9),
    502 => to_signed(0, 9),
    503 => to_signed(8, 9),
    504 => to_signed(-2, 9),
    505 => to_signed(-16, 9),
    506 => to_signed(5, 9),
    507 => to_signed(19, 9),
    508 => to_signed(-7, 9),
    509 => to_signed(1, 9),
    510 => to_signed(4, 9),
    511 => to_signed(1, 9),
    512 => to_signed(4, 9),
    513 => to_signed(51, 9),
    514 => to_signed(32, 9),
    515 => to_signed(21, 9),
    516 => to_signed(3, 9),
    517 => to_signed(2, 9),
    518 => to_signed(0, 9),
    519 => to_signed(0, 9),
    520 => to_signed(26, 9),
    521 => to_signed(56, 9),
    522 => to_signed(43, 9),
    523 => to_signed(18, 9),
    524 => to_signed(-10, 9),
    525 => to_signed(2, 9),
    526 => to_signed(0, 9),
    527 => to_signed(1, 9),
    528 => to_signed(16, 9),
    529 => to_signed(57, 9),
    530 => to_signed(14, 9),
    531 => to_signed(25, 9),
    532 => to_signed(0, 9),
    533 => to_signed(-2, 9),
    534 => to_signed(2, 9),
    535 => to_signed(11, 9),
    536 => to_signed(-52, 9),
    537 => to_signed(-48, 9),
    538 => to_signed(28, 9),
    539 => to_signed(26, 9),
    540 => to_signed(31, 9),
    541 => to_signed(-4, 9),
    542 => to_signed(-5, 9),
    543 => to_signed(1, 9),
    544 => to_signed(-1, 9),
    545 => to_signed(-55, 9),
    546 => to_signed(-52, 9),
    547 => to_signed(-18, 9),
    548 => to_signed(5, 9),
    549 => to_signed(-5, 9),
    550 => to_signed(0, 9),
    551 => to_signed(0, 9),
    552 => to_signed(-2, 9),
    553 => to_signed(4, 9),
    554 => to_signed(-3, 9),
    555 => to_signed(-39, 9),
    556 => to_signed(-59, 9),
    557 => to_signed(-19, 9),
    558 => to_signed(0, 9),
    559 => to_signed(-1, 9),
    560 => to_signed(-3, 9),
    561 => to_signed(0, 9),
    562 => to_signed(-3, 9),
    563 => to_signed(1, 9),
    564 => to_signed(2, 9),
    565 => to_signed(-2, 9),
    566 => to_signed(2, 9),
    567 => to_signed(0, 9),
    568 => to_signed(-4, 9),
    569 => to_signed(0, 9),
    570 => to_signed(0, 9),
    571 => to_signed(1, 9),
    572 => to_signed(0, 9),
    573 => to_signed(1, 9),
    574 => to_signed(1, 9),
    575 => to_signed(-2, 9),
    576 => to_signed(0, 9),
    577 => to_signed(-2, 9),
    578 => to_signed(0, 9),
    579 => to_signed(-2, 9),
    580 => to_signed(-1, 9),
    581 => to_signed(0, 9),
    582 => to_signed(-1, 9),
    583 => to_signed(-1, 9),
    584 => to_signed(1, 9),
    585 => to_signed(-2, 9),
    586 => to_signed(3, 9),
    587 => to_signed(-1, 9),
    588 => to_signed(-4, 9),
    589 => to_signed(0, 9),
    590 => to_signed(2, 9),
    591 => to_signed(-6, 9),
    592 => to_signed(1, 9),
    593 => to_signed(-5, 9),
    594 => to_signed(-4, 9),
    595 => to_signed(-3, 9),
    596 => to_signed(-3, 9),
    597 => to_signed(1, 9),
    598 => to_signed(1, 9),
    599 => to_signed(0, 9),
    600 => to_signed(4, 9),
    601 => to_signed(2, 9),
    602 => to_signed(-4, 9),
    603 => to_signed(-7, 9),
    604 => to_signed(0, 9),
    605 => to_signed(-1, 9),
    606 => to_signed(2, 9),
    607 => to_signed(0, 9),
    608 => to_signed(0, 9),
    609 => to_signed(0, 9),
    610 => to_signed(-1, 9),
    611 => to_signed(0, 9),
    612 => to_signed(0, 9),
    613 => to_signed(0, 9),
    614 => to_signed(-2, 9),
    615 => to_signed(0, 9),
    616 => to_signed(-3, 9),
    617 => to_signed(0, 9),
    618 => to_signed(0, 9),
    619 => to_signed(0, 9),
    620 => to_signed(0, 9),
    621 => to_signed(1, 9),
    622 => to_signed(4, 9),
    623 => to_signed(0, 9),
    624 => to_signed(-3, 9),
    625 => to_signed(0, 9),
    626 => to_signed(0, 9),
    627 => to_signed(-1, 9),
    628 => to_signed(0, 9),
    629 => to_signed(1, 9),
    630 => to_signed(-3, 9),
    631 => to_signed(0, 9),
    632 => to_signed(-2, 9),
    633 => to_signed(5, 9),
    634 => to_signed(2, 9),
    635 => to_signed(-2, 9),
    636 => to_signed(0, 9),
    637 => to_signed(0, 9),
    638 => to_signed(0, 9),
    639 => to_signed(0, 9),
    640 => to_signed(0, 9),
    641 => to_signed(-1, 9),
    642 => to_signed(6, 9),
    643 => to_signed(5, 9),
    644 => to_signed(2, 9),
    645 => to_signed(0, 9),
    646 => to_signed(-6, 9),
    647 => to_signed(-1, 9),
    648 => to_signed(1, 9),
    649 => to_signed(0, 9),
    650 => to_signed(0, 9),
    651 => to_signed(-2, 9),
    652 => to_signed(-3, 9),
    653 => to_signed(-4, 9),
    654 => to_signed(0, 9),
    655 => to_signed(-4, 9),
    656 => to_signed(0, 9),
    657 => to_signed(-1, 9),
    658 => to_signed(-1, 9),
    659 => to_signed(-3, 9),
    660 => to_signed(-2, 9),
    661 => to_signed(1, 9),
    662 => to_signed(-1, 9),
    663 => to_signed(0, 9),
    664 => to_signed(-1, 9),
    665 => to_signed(0, 9),
    666 => to_signed(0, 9),
    667 => to_signed(-1, 9),
    668 => to_signed(1, 9),
    669 => to_signed(0, 9),
    670 => to_signed(-3, 9),
    671 => to_signed(-1, 9),
    672 => to_signed(0, 9),
    673 => to_signed(-1, 9),
    674 => to_signed(-6, 9),
    675 => to_signed(-3, 9),
    676 => to_signed(-6, 9),
    677 => to_signed(-2, 9),
    678 => to_signed(2, 9),
    679 => to_signed(0, 9),
    680 => to_signed(2, 9),
    681 => to_signed(-2, 9),
    682 => to_signed(8, 9),
    683 => to_signed(0, 9),
    684 => to_signed(3, 9),
    685 => to_signed(7, 9),
    686 => to_signed(5, 9),
    687 => to_signed(1, 9),
    688 => to_signed(-3, 9),
    689 => to_signed(10, 9),
    690 => to_signed(14, 9),
    691 => to_signed(9, 9),
    692 => to_signed(2, 9),
    693 => to_signed(3, 9),
    694 => to_signed(-4, 9),
    695 => to_signed(3, 9),
    696 => to_signed(1, 9),
    697 => to_signed(7, 9),
    698 => to_signed(-12, 9),
    699 => to_signed(-31, 9),
    700 => to_signed(-9, 9),
    701 => to_signed(6, 9),
    702 => to_signed(8, 9),
    703 => to_signed(-1, 9),
    704 => to_signed(-1, 9),
    705 => to_signed(-11, 9),
    706 => to_signed(-21, 9),
    707 => to_signed(0, 9),
    708 => to_signed(1, 9),
    709 => to_signed(-4, 9),
    710 => to_signed(1, 9),
    711 => to_signed(-4, 9),
    712 => to_signed(0, 9),
    713 => to_signed(-6, 9),
    714 => to_signed(-4, 9),
    715 => to_signed(15, 9),
    716 => to_signed(1, 9),
    717 => to_signed(-13, 9),
    718 => to_signed(-6, 9),
    719 => to_signed(-2, 9),
    720 => to_signed(2, 9),
    721 => to_signed(1, 9),
    722 => to_signed(21, 9),
    723 => to_signed(10, 9),
    724 => to_signed(1, 9),
    725 => to_signed(-3, 9),
    726 => to_signed(-2, 9),
    727 => to_signed(5, 9),
    728 => to_signed(-2, 9),
    729 => to_signed(6, 9),
    730 => to_signed(11, 9),
    731 => to_signed(-1, 9),
    732 => to_signed(12, 9),
    733 => to_signed(10, 9),
    734 => to_signed(-4, 9),
    735 => to_signed(-3, 9),
    736 => to_signed(-2, 9),
    737 => to_signed(3, 9),
    738 => to_signed(12, 9),
    739 => to_signed(13, 9),
    740 => to_signed(2, 9),
    741 => to_signed(-8, 9),
    742 => to_signed(2, 9),
    743 => to_signed(1, 9),
    744 => to_signed(2, 9),
    745 => to_signed(6, 9),
    746 => to_signed(-20, 9),
    747 => to_signed(-29, 9),
    748 => to_signed(-12, 9),
    749 => to_signed(-4, 9),
    750 => to_signed(-2, 9),
    751 => to_signed(4, 9),
    752 => to_signed(7, 9),
    753 => to_signed(6, 9),
    754 => to_signed(18, 9),
    755 => to_signed(-7, 9),
    756 => to_signed(3, 9),
    757 => to_signed(1, 9),
    758 => to_signed(2, 9),
    759 => to_signed(3, 9),
    760 => to_signed(-7, 9),
    761 => to_signed(-2, 9),
    762 => to_signed(13, 9),
    763 => to_signed(27, 9),
    764 => to_signed(17, 9),
    765 => to_signed(-4, 9),
    766 => to_signed(0, 9),
    767 => to_signed(6, 9),
    768 => to_signed(-16, 9),
    769 => to_signed(-31, 9),
    770 => to_signed(-22, 9),
    771 => to_signed(-4, 9),
    772 => to_signed(1, 9),
    773 => to_signed(1, 9),
    774 => to_signed(-3, 9),
    775 => to_signed(3, 9),
    776 => to_signed(-1, 9),
    777 => to_signed(-39, 9),
    778 => to_signed(-3, 9),
    779 => to_signed(-7, 9),
    780 => to_signed(-8, 9),
    781 => to_signed(0, 9),
    782 => to_signed(-2, 9),
    783 => to_signed(2, 9),
    784 => to_signed(42, 9),
    785 => to_signed(16, 9),
    786 => to_signed(-6, 9),
    787 => to_signed(8, 9),
    788 => to_signed(-15, 9),
    789 => to_signed(0, 9),
    790 => to_signed(-2, 9),
    791 => to_signed(4, 9),
    792 => to_signed(18, 9),
    793 => to_signed(40, 9),
    794 => to_signed(48, 9),
    795 => to_signed(37, 9),
    796 => to_signed(-15, 9),
    797 => to_signed(2, 9),
    798 => to_signed(-1, 9),
    799 => to_signed(11, 9),
    800 => to_signed(12, 9),
    801 => to_signed(11, 9),
    802 => to_signed(13, 9),
    803 => to_signed(12, 9),
    804 => to_signed(14, 9),
    805 => to_signed(5, 9),
    806 => to_signed(0, 9),
    807 => to_signed(2, 9),
    808 => to_signed(10, 9),
    809 => to_signed(3, 9),
    810 => to_signed(0, 9),
    811 => to_signed(-3, 9),
    812 => to_signed(3, 9),
    813 => to_signed(16, 9),
    814 => to_signed(12, 9),
    815 => to_signed(3, 9),
    816 => to_signed(1, 9),
    817 => to_signed(5, 9),
    818 => to_signed(7, 9),
    819 => to_signed(-1, 9),
    820 => to_signed(-4, 9),
    821 => to_signed(1, 9),
    822 => to_signed(-31, 9),
    823 => to_signed(-26, 9),
    824 => to_signed(-1, 9),
    825 => to_signed(1, 9),
    826 => to_signed(8, 9),
    827 => to_signed(2, 9),
    828 => to_signed(1, 9),
    829 => to_signed(-6, 9),
    830 => to_signed(-29, 9),
    831 => to_signed(3, 9),
    832 => to_signed(14, 9),
    833 => to_signed(-22, 9),
    834 => to_signed(-9, 9),
    835 => to_signed(-2, 9),
    836 => to_signed(-1, 9),
    837 => to_signed(-2, 9),
    838 => to_signed(-8, 9),
    839 => to_signed(16, 9),
    840 => to_signed(19, 9),
    841 => to_signed(6, 9),
    842 => to_signed(-1, 9),
    843 => to_signed(-2, 9),
    844 => to_signed(-2, 9),
    845 => to_signed(-7, 9),
    846 => to_signed(-5, 9),
    847 => to_signed(-15, 9),
    848 => to_signed(9, 9),
    849 => to_signed(19, 9),
    850 => to_signed(12, 9),
    851 => to_signed(-1, 9),
    852 => to_signed(-2, 9),
    853 => to_signed(0, 9),
    854 => to_signed(11, 9),
    855 => to_signed(4, 9),
    856 => to_signed(17, 9),
    857 => to_signed(30, 9),
    858 => to_signed(-6, 9),
    859 => to_signed(-1, 9),
    860 => to_signed(-1, 9),
    861 => to_signed(11, 9),
    862 => to_signed(17, 9),
    863 => to_signed(12, 9),
    864 => to_signed(0, 9),
    865 => to_signed(-5, 9),
    866 => to_signed(-14, 9),
    867 => to_signed(-5, 9),
    868 => to_signed(-4, 9),
    869 => to_signed(7, 9),
    870 => to_signed(-13, 9),
    871 => to_signed(-10, 9),
    872 => to_signed(5, 9),
    873 => to_signed(3, 9),
    874 => to_signed(1, 9),
    875 => to_signed(-24, 9),
    876 => to_signed(-6, 9),
    877 => to_signed(-11, 9),
    878 => to_signed(-42, 9),
    879 => to_signed(-15, 9),
    880 => to_signed(9, 9),
    881 => to_signed(0, 9),
    882 => to_signed(1, 9),
    883 => to_signed(-22, 9),
    884 => to_signed(11, 9),
    885 => to_signed(-10, 9),
    886 => to_signed(-14, 9),
    887 => to_signed(-50, 9),
    888 => to_signed(-6, 9),
    889 => to_signed(0, 9),
    890 => to_signed(0, 9),
    891 => to_signed(-15, 9),
    892 => to_signed(7, 9),
    893 => to_signed(0, 9),
    894 => to_signed(28, 9),
    895 => to_signed(-34, 9),
    896 => to_signed(-25, 9),
    897 => to_signed(0, 9),
    898 => to_signed(-2, 9),
    899 => to_signed(1, 9),
    900 => to_signed(18, 9),
    901 => to_signed(34, 9),
    902 => to_signed(25, 9),
    903 => to_signed(-2, 9),
    904 => to_signed(-12, 9),
    905 => to_signed(2, 9),
    906 => to_signed(0, 9),
    907 => to_signed(-13, 9),
    908 => to_signed(81, 9),
    909 => to_signed(89, 9),
    910 => to_signed(-4, 9),
    911 => to_signed(-25, 9),
    912 => to_signed(10, 9),
    913 => to_signed(1, 9),
    914 => to_signed(1, 9),
    915 => to_signed(-30, 9),
    916 => to_signed(28, 9),
    917 => to_signed(39, 9),
    918 => to_signed(-16, 9),
    919 => to_signed(-9, 9),
    920 => to_signed(6, 9),
    921 => to_signed(7, 9),
    922 => to_signed(-4, 9),
    923 => to_signed(-5, 9),
    924 => to_signed(-3, 9),
    925 => to_signed(5, 9),
    926 => to_signed(-1, 9),
    927 => to_signed(26, 9),
    928 => to_signed(16, 9),
    929 => to_signed(7, 9),
    930 => to_signed(3, 9),
    931 => to_signed(1, 9),
    932 => to_signed(26, 9),
    933 => to_signed(19, 9),
    934 => to_signed(16, 9),
    935 => to_signed(-5, 9),
    936 => to_signed(0, 9),
    937 => to_signed(3, 9),
    938 => to_signed(5, 9),
    939 => to_signed(0, 9),
    940 => to_signed(-16, 9),
    941 => to_signed(11, 9),
    942 => to_signed(14, 9),
    943 => to_signed(0, 9),
    944 => to_signed(0, 9),
    945 => to_signed(-8, 9),
    946 => to_signed(-18, 9),
    947 => to_signed(0, 9),
    948 => to_signed(2, 9),
    949 => to_signed(-21, 9),
    950 => to_signed(-7, 9),
    951 => to_signed(4, 9),
    952 => to_signed(-2, 9),
    953 => to_signed(-9, 9),
    954 => to_signed(-7, 9),
    955 => to_signed(16, 9),
    956 => to_signed(30, 9),
    957 => to_signed(-20, 9),
    958 => to_signed(-34, 9),
    959 => to_signed(2, 9),
    960 => to_signed(1, 9),
    961 => to_signed(-5, 9),
    962 => to_signed(-21, 9),
    963 => to_signed(14, 9),
    964 => to_signed(8, 9),
    965 => to_signed(10, 9),
    966 => to_signed(-8, 9),
    967 => to_signed(-1, 9),
    968 => to_signed(1, 9),
    969 => to_signed(-28, 9),
    970 => to_signed(-66, 9),
    971 => to_signed(-38, 9),
    972 => to_signed(-10, 9),
    973 => to_signed(16, 9),
    974 => to_signed(39, 9),
    975 => to_signed(2, 9),
    976 => to_signed(0, 9),
    977 => to_signed(-17, 9),
    978 => to_signed(-4, 9),
    979 => to_signed(-1, 9),
    980 => to_signed(-5, 9),
    981 => to_signed(36, 9),
    982 => to_signed(28, 9),
    983 => to_signed(1, 9),
    984 => to_signed(-2, 9),
    985 => to_signed(10, 9),
    986 => to_signed(22, 9),
    987 => to_signed(29, 9),
    988 => to_signed(24, 9),
    989 => to_signed(27, 9),
    990 => to_signed(0, 9),
    991 => to_signed(-3, 9),
    992 => to_signed(-4, 9),
    993 => to_signed(0, 9),
    994 => to_signed(7, 9),
    995 => to_signed(-4, 9),
    996 => to_signed(-4, 9),
    997 => to_signed(0, 9),
    998 => to_signed(-2, 9),
    999 => to_signed(-3, 9),
    1000 => to_signed(-3, 9),
    1001 => to_signed(1, 9),
    1002 => to_signed(3, 9),
    1003 => to_signed(4, 9),
    1004 => to_signed(-3, 9),
    1005 => to_signed(1, 9),
    1006 => to_signed(1, 9),
    1007 => to_signed(-2, 9),
    1008 => to_signed(2, 9),
    1009 => to_signed(-2, 9),
    1010 => to_signed(0, 9),
    1011 => to_signed(-5, 9),
    1012 => to_signed(0, 9),
    1013 => to_signed(-6, 9),
    1014 => to_signed(0, 9),
    1015 => to_signed(0, 9),
    1016 => to_signed(4, 9),
    1017 => to_signed(-2, 9),
    1018 => to_signed(1, 9),
    1019 => to_signed(-1, 9),
    1020 => to_signed(1, 9),
    1021 => to_signed(-1, 9),
    1022 => to_signed(3, 9),
    1023 => to_signed(0, 9),
    1024 => to_signed(3, 9),
    1025 => to_signed(5, 9),
    1026 => to_signed(-2, 9),
    1027 => to_signed(6, 9),
    1028 => to_signed(-2, 9),
    1029 => to_signed(0, 9),
    1030 => to_signed(5, 9),
    1031 => to_signed(-4, 9),
    1032 => to_signed(4, 9),
    1033 => to_signed(4, 9),
    1034 => to_signed(-5, 9),
    1035 => to_signed(-2, 9),
    1036 => to_signed(4, 9),
    1037 => to_signed(1, 9),
    1038 => to_signed(0, 9),
    1039 => to_signed(-7, 9),
    1040 => to_signed(-4, 9),
    1041 => to_signed(-1, 9),
    1042 => to_signed(-1, 9),
    1043 => to_signed(-4, 9),
    1044 => to_signed(3, 9),
    1045 => to_signed(0, 9),
    1046 => to_signed(0, 9),
    1047 => to_signed(2, 9),
    1048 => to_signed(-2, 9),
    1049 => to_signed(0, 9),
    1050 => to_signed(1, 9),
    1051 => to_signed(5, 9),
    1052 => to_signed(4, 9),
    1053 => to_signed(-1, 9),
    1054 => to_signed(10, 9),
    1055 => to_signed(9, 9),
    1056 => to_signed(17, 9),
    1057 => to_signed(-17, 9),
    1058 => to_signed(-12, 9),
    1059 => to_signed(-8, 9),
    1060 => to_signed(-1, 9),
    1061 => to_signed(14, 9),
    1062 => to_signed(16, 9),
    1063 => to_signed(-17, 9),
    1064 => to_signed(12, 9),
    1065 => to_signed(13, 9),
    1066 => to_signed(21, 9),
    1067 => to_signed(3, 9),
    1068 => to_signed(0, 9),
    1069 => to_signed(8, 9),
    1070 => to_signed(-34, 9),
    1071 => to_signed(-28, 9),
    1072 => to_signed(46, 9),
    1073 => to_signed(47, 9),
    1074 => to_signed(29, 9),
    1075 => to_signed(3, 9),
    1076 => to_signed(-2, 9),
    1077 => to_signed(-6, 9),
    1078 => to_signed(-35, 9),
    1079 => to_signed(-11, 9),
    1080 => to_signed(39, 9),
    1081 => to_signed(32, 9),
    1082 => to_signed(16, 9),
    1083 => to_signed(-1, 9),
    1084 => to_signed(-2, 9),
    1085 => to_signed(-9, 9),
    1086 => to_signed(-19, 9),
    1087 => to_signed(-1, 9),
    1088 => to_signed(51, 9),
    1089 => to_signed(52, 9),
    1090 => to_signed(0, 9),
    1091 => to_signed(1, 9),
    1092 => to_signed(1, 9),
    1093 => to_signed(7, 9),
    1094 => to_signed(-53, 9),
    1095 => to_signed(-6, 9),
    1096 => to_signed(26, 9),
    1097 => to_signed(-8, 9),
    1098 => to_signed(-19, 9),
    1099 => to_signed(-5, 9),
    1100 => to_signed(-2, 9),
    1101 => to_signed(9, 9),
    1102 => to_signed(-35, 9),
    1103 => to_signed(-26, 9),
    1104 => to_signed(-24, 9),
    1105 => to_signed(-5, 9),
    1106 => to_signed(-3, 9),
    1107 => to_signed(-3, 9),
    1108 => to_signed(0, 9),
    1109 => to_signed(2, 9),
    1110 => to_signed(12, 9),
    1111 => to_signed(-21, 9),
    1112 => to_signed(-2, 9),
    1113 => to_signed(26, 9),
    1114 => to_signed(1, 9),
    1115 => to_signed(8, 9),
    1116 => to_signed(6, 9),
    1117 => to_signed(-7, 9),
    1118 => to_signed(-13, 9),
    1119 => to_signed(-12, 9),
    1120 => to_signed(-1, 9),
    1121 => to_signed(0, 9),
    1122 => to_signed(-4, 9),
    1123 => to_signed(-8, 9),
    1124 => to_signed(-18, 9),
    1125 => to_signed(-15, 9),
    1126 => to_signed(-43, 9),
    1127 => to_signed(-31, 9),
    1128 => to_signed(14, 9),
    1129 => to_signed(1, 9),
    1130 => to_signed(3, 9),
    1131 => to_signed(-2, 9),
    1132 => to_signed(10, 9),
    1133 => to_signed(15, 9),
    1134 => to_signed(2, 9),
    1135 => to_signed(-44, 9),
    1136 => to_signed(0, 9),
    1137 => to_signed(-1, 9),
    1138 => to_signed(0, 9),
    1139 => to_signed(0, 9),
    1140 => to_signed(4, 9),
    1141 => to_signed(8, 9),
    1142 => to_signed(17, 9),
    1143 => to_signed(-21, 9),
    1144 => to_signed(-14, 9),
    1145 => to_signed(0, 9),
    1146 => to_signed(0, 9),
    1147 => to_signed(8, 9),
    1148 => to_signed(1, 9),
    1149 => to_signed(-9, 9),
    1150 => to_signed(21, 9),
    1151 => to_signed(9, 9),
    1152 => to_signed(-7, 9),
    1153 => to_signed(1, 9),
    1154 => to_signed(1, 9),
    1155 => to_signed(-5, 9),
    1156 => to_signed(19, 9),
    1157 => to_signed(46, 9),
    1158 => to_signed(20, 9),
    1159 => to_signed(-4, 9),
    1160 => to_signed(-6, 9),
    1161 => to_signed(-2, 9),
    1162 => to_signed(1, 9),
    1163 => to_signed(-2, 9),
    1164 => to_signed(1, 9),
    1165 => to_signed(34, 9),
    1166 => to_signed(22, 9),
    1167 => to_signed(18, 9),
    1168 => to_signed(18, 9),
    1169 => to_signed(7, 9),
    1170 => to_signed(1, 9),
    1171 => to_signed(0, 9),
    1172 => to_signed(15, 9),
    1173 => to_signed(-1, 9),
    1174 => to_signed(10, 9),
    1175 => to_signed(49, 9),
    1176 => to_signed(37, 9),
    1177 => to_signed(8, 9),
    1178 => to_signed(7, 9),
    1179 => to_signed(17, 9),
    1180 => to_signed(21, 9),
    1181 => to_signed(17, 9),
    1182 => to_signed(6, 9),
    1183 => to_signed(3, 9),
    1184 => to_signed(3, 9),
    1185 => to_signed(11, 9),
    1186 => to_signed(29, 9),
    1187 => to_signed(20, 9),
    1188 => to_signed(8, 9),
    1189 => to_signed(12, 9),
    1190 => to_signed(2, 9),
    1191 => to_signed(6, 9),
    1192 => to_signed(0, 9),
    1193 => to_signed(-2, 9),
    1194 => to_signed(-5, 9),
    1195 => to_signed(-42, 9),
    1196 => to_signed(-13, 9),
    1197 => to_signed(22, 9),
    1198 => to_signed(13, 9),
    1199 => to_signed(1, 9),
    1200 => to_signed(-1, 9),
    1201 => to_signed(-10, 9),
    1202 => to_signed(-11, 9),
    1203 => to_signed(0, 9),
    1204 => to_signed(15, 9),
    1205 => to_signed(19, 9),
    1206 => to_signed(17, 9),
    1207 => to_signed(-4, 9),
    1208 => to_signed(0, 9),
    1209 => to_signed(0, 9),
    1210 => to_signed(0, 9),
    1211 => to_signed(23, 9),
    1212 => to_signed(12, 9),
    1213 => to_signed(3, 9),
    1214 => to_signed(5, 9),
    1215 => to_signed(3, 9),
    1216 => to_signed(5, 9),
    1217 => to_signed(6, 9),
    1218 => to_signed(8, 9),
    1219 => to_signed(-2, 9),
    1220 => to_signed(-2, 9),
    1221 => to_signed(-9, 9),
    1222 => to_signed(2, 9),
    1223 => to_signed(0, 9),
    1224 => to_signed(-3, 9),
    1225 => to_signed(3, 9),
    1226 => to_signed(-3, 9),
    1227 => to_signed(-17, 9),
    1228 => to_signed(-38, 9),
    1229 => to_signed(-25, 9),
    1230 => to_signed(6, 9),
    1231 => to_signed(4, 9),
    1232 => to_signed(0, 9),
    1233 => to_signed(-2, 9),
    1234 => to_signed(0, 9),
    1235 => to_signed(2, 9),
    1236 => to_signed(-16, 9),
    1237 => to_signed(-22, 9),
    1238 => to_signed(1, 9),
    1239 => to_signed(-2, 9),
    1240 => to_signed(-27, 9),
    1241 => to_signed(29, 9),
    1242 => to_signed(7, 9),
    1243 => to_signed(6, 9),
    1244 => to_signed(-11, 9),
    1245 => to_signed(-12, 9),
    1246 => to_signed(5, 9),
    1247 => to_signed(22, 9),
    1248 => to_signed(26, 9),
    1249 => to_signed(1, 9),
    1250 => to_signed(17, 9),
    1251 => to_signed(29, 9),
    1252 => to_signed(-13, 9),
    1253 => to_signed(2, 9),
    1254 => to_signed(1, 9),
    1255 => to_signed(4, 9),
    1256 => to_signed(-4, 9),
    1257 => to_signed(-45, 9),
    1258 => to_signed(0, 9),
    1259 => to_signed(55, 9),
    1260 => to_signed(36, 9),
    1261 => to_signed(0, 9),
    1262 => to_signed(-2, 9),
    1263 => to_signed(-24, 9),
    1264 => to_signed(-25, 9),
    1265 => to_signed(-26, 9),
    1266 => to_signed(15, 9),
    1267 => to_signed(20, 9),
    1268 => to_signed(-4, 9),
    1269 => to_signed(2, 9),
    1270 => to_signed(0, 9),
    1271 => to_signed(-19, 9),
    1272 => to_signed(7, 9),
    1273 => to_signed(35, 9),
    1274 => to_signed(8, 9),
    1275 => to_signed(-5, 9),
    1276 => to_signed(-33, 9),
    1277 => to_signed(1, 9),
    1278 => to_signed(2, 9),
    1279 => to_signed(-13, 9),
    1280 => to_signed(72, 9),
    1281 => to_signed(19, 9),
    1282 => to_signed(-12, 9),
    1283 => to_signed(-7, 9),
    1284 => to_signed(-18, 9),
    1285 => to_signed(-1, 9),
    1286 => to_signed(-2, 9),
    1287 => to_signed(-16, 9),
    1288 => to_signed(8, 9),
    1289 => to_signed(-15, 9),
    1290 => to_signed(-22, 9),
    1291 => to_signed(-3, 9),
    1292 => to_signed(-2, 9),
    1293 => to_signed(0, 9),
    1294 => to_signed(1, 9),
    1295 => to_signed(0, 9),
    1296 => to_signed(-20, 9),
    1297 => to_signed(27, 9),
    1298 => to_signed(6, 9),
    1299 => to_signed(10, 9),
    1300 => to_signed(28, 9),
    1301 => to_signed(0, 9),
    1302 => to_signed(19, 9),
    1303 => to_signed(9, 9),
    1304 => to_signed(25, 9),
    1305 => to_signed(4, 9),
    1306 => to_signed(-12, 9),
    1307 => to_signed(-2, 9),
    1308 => to_signed(-1, 9),
    1309 => to_signed(10, 9),
    1310 => to_signed(13, 9),
    1311 => to_signed(0, 9),
    1312 => to_signed(25, 9),
    1313 => to_signed(13, 9),
    1314 => to_signed(0, 9),
    1315 => to_signed(0, 9),
    1316 => to_signed(-2, 9),
    1317 => to_signed(-20, 9),
    1318 => to_signed(-65, 9),
    1319 => to_signed(-57, 9),
    1320 => to_signed(43, 9),
    1321 => to_signed(13, 9),
    1322 => to_signed(2, 9),
    1323 => to_signed(6, 9),
    1324 => to_signed(1, 9),
    1325 => to_signed(-12, 9),
    1326 => to_signed(-43, 9),
    1327 => to_signed(2, 9),
    1328 => to_signed(38, 9),
    1329 => to_signed(13, 9),
    1330 => to_signed(28, 9),
    1331 => to_signed(1, 9),
    1332 => to_signed(-2, 9),
    1333 => to_signed(0, 9),
    1334 => to_signed(18, 9),
    1335 => to_signed(20, 9),
    1336 => to_signed(50, 9),
    1337 => to_signed(18, 9),
    1338 => to_signed(13, 9),
    1339 => to_signed(4, 9),
    1340 => to_signed(-1, 9),
    1341 => to_signed(24, 9),
    1342 => to_signed(12, 9),
    1343 => to_signed(34, 9),
    1344 => to_signed(20, 9),
    1345 => to_signed(-35, 9),
    1346 => to_signed(-21, 9),
    1347 => to_signed(1, 9),
    1348 => to_signed(0, 9),
    1349 => to_signed(36, 9),
    1350 => to_signed(12, 9),
    1351 => to_signed(-3, 9),
    1352 => to_signed(-27, 9),
    1353 => to_signed(-21, 9),
    1354 => to_signed(-22, 9),
    1355 => to_signed(-8, 9),
    1356 => to_signed(-4, 9),
    1357 => to_signed(4, 9),
    1358 => to_signed(18, 9),
    1359 => to_signed(-24, 9),
    1360 => to_signed(-38, 9),
    1361 => to_signed(-17, 9),
    1362 => to_signed(-10, 9),
    1363 => to_signed(7, 9),
    1364 => to_signed(-23, 9),
    1365 => to_signed(-7, 9),
    1366 => to_signed(4, 9),
    1367 => to_signed(7, 9),
    1368 => to_signed(-13, 9),
    1369 => to_signed(3, 9),
    1370 => to_signed(4, 9),
    1371 => to_signed(0, 9),
    1372 => to_signed(8, 9),
    1373 => to_signed(0, 9),
    1374 => to_signed(-15, 9),
    1375 => to_signed(14, 9),
    1376 => to_signed(-10, 9),
    1377 => to_signed(-2, 9),
    1378 => to_signed(-2, 9),
    1379 => to_signed(21, 9),
    1380 => to_signed(28, 9),
    1381 => to_signed(-29, 9),
    1382 => to_signed(-38, 9),
    1383 => to_signed(2, 9),
    1384 => to_signed(0, 9),
    1385 => to_signed(0, 9),
    1386 => to_signed(3, 9),
    1387 => to_signed(1, 9),
    1388 => to_signed(-8, 9),
    1389 => to_signed(-23, 9),
    1390 => to_signed(-20, 9),
    1391 => to_signed(-19, 9),
    1392 => to_signed(-16, 9),
    1393 => to_signed(0, 9),
    1394 => to_signed(0, 9),
    1395 => to_signed(-4, 9),
    1396 => to_signed(0, 9),
    1397 => to_signed(-1, 9),
    1398 => to_signed(-14, 9),
    1399 => to_signed(-35, 9),
    1400 => to_signed(-15, 9),
    1401 => to_signed(2, 9),
    1402 => to_signed(1, 9),
    1403 => to_signed(-12, 9),
    1404 => to_signed(84, 9),
    1405 => to_signed(27, 9),
    1406 => to_signed(-7, 9),
    1407 => to_signed(0, 9),
    1408 => to_signed(11, 9),
    1409 => to_signed(2, 9),
    1410 => to_signed(-3, 9),
    1411 => to_signed(-23, 9),
    1412 => to_signed(30, 9),
    1413 => to_signed(14, 9),
    1414 => to_signed(27, 9),
    1415 => to_signed(38, 9),
    1416 => to_signed(12, 9),
    1417 => to_signed(6, 9),
    1418 => to_signed(2, 9),
    1419 => to_signed(2, 9),
    1420 => to_signed(-13, 9),
    1421 => to_signed(25, 9),
    1422 => to_signed(32, 9),
    1423 => to_signed(21, 9),
    1424 => to_signed(20, 9),
    1425 => to_signed(3, 9),
    1426 => to_signed(5, 9),
    1427 => to_signed(5, 9),
    1428 => to_signed(1, 9),
    1429 => to_signed(0, 9),
    1430 => to_signed(2, 9),
    1431 => to_signed(1, 9),
    1432 => to_signed(0, 9),
    1433 => to_signed(3, 9),
    1434 => to_signed(1, 9),
    1435 => to_signed(13, 9),
    1436 => to_signed(15, 9),
    1437 => to_signed(-3, 9),
    1438 => to_signed(-2, 9),
    1439 => to_signed(0, 9),
    1440 => to_signed(-1, 9),
    1441 => to_signed(0, 9),
    1442 => to_signed(1, 9),
    1443 => to_signed(16, 9),
    1444 => to_signed(14, 9),
    1445 => to_signed(-14, 9),
    1446 => to_signed(-6, 9),
    1447 => to_signed(-3, 9),
    1448 => to_signed(-1, 9),
    1449 => to_signed(-2, 9),
    1450 => to_signed(-2, 9),
    1451 => to_signed(-7, 9),
    1452 => to_signed(0, 9),
    1453 => to_signed(-5, 9),
    1454 => to_signed(-8, 9),
    1455 => to_signed(-3, 9),
    1456 => to_signed(1, 9),
    1457 => to_signed(-1, 9),
    1458 => to_signed(-6, 9),
    1459 => to_signed(-2, 9),
    1460 => to_signed(-4, 9),
    1461 => to_signed(-4, 9),
    1462 => to_signed(2, 9),
    1463 => to_signed(-2, 9),
    1464 => to_signed(-3, 9),
    1465 => to_signed(-13, 9),
    1466 => to_signed(-14, 9),
    1467 => to_signed(2, 9),
    1468 => to_signed(-4, 9),
    1469 => to_signed(-14, 9),
    1470 => to_signed(-5, 9),
    1471 => to_signed(0, 9),
    1472 => to_signed(1, 9),
    1473 => to_signed(-11, 9),
    1474 => to_signed(-10, 9),
    1475 => to_signed(4, 9),
    1476 => to_signed(10, 9),
    1477 => to_signed(-2, 9),
    1478 => to_signed(-2, 9),
    1479 => to_signed(1, 9),
    1480 => to_signed(-3, 9),
    1481 => to_signed(3, 9),
    1482 => to_signed(3, 9),
    1483 => to_signed(4, 9),
    1484 => to_signed(6, 9),
    1485 => to_signed(17, 9),
    1486 => to_signed(7, 9),
    1487 => to_signed(-3, 9),
    1488 => to_signed(3, 9),
    1489 => to_signed(-2, 9),
    1490 => to_signed(-33, 9),
    1491 => to_signed(-10, 9),
    1492 => to_signed(-3, 9),
    1493 => to_signed(1, 9),
    1494 => to_signed(-5, 9),
    1495 => to_signed(-34, 9),
    1496 => to_signed(-40, 9),
    1497 => to_signed(-19, 9),
    1498 => to_signed(-2, 9),
    1499 => to_signed(6, 9),
    1500 => to_signed(10, 9),
    1501 => to_signed(-8, 9),
    1502 => to_signed(1, 9),
    1503 => to_signed(5, 9),
    1504 => to_signed(47, 9),
    1505 => to_signed(105, 9),
    1506 => to_signed(54, 9),
    1507 => to_signed(39, 9),
    1508 => to_signed(-4, 9),
    1509 => to_signed(-4, 9),
    1510 => to_signed(-2, 9),
    1511 => to_signed(7, 9),
    1512 => to_signed(52, 9),
    1513 => to_signed(12, 9),
    1514 => to_signed(-1, 9),
    1515 => to_signed(62, 9),
    1516 => to_signed(6, 9),
    1517 => to_signed(1, 9),
    1518 => to_signed(-5, 9),
    1519 => to_signed(6, 9),
    1520 => to_signed(13, 9),
    1521 => to_signed(-26, 9),
    1522 => to_signed(-15, 9),
    1523 => to_signed(10, 9),
    1524 => to_signed(0, 9),
    1525 => to_signed(-3, 9),
    1526 => to_signed(0, 9),
    1527 => to_signed(16, 9),
    1528 => to_signed(-32, 9),
    1529 => to_signed(8, 9),
    1530 => to_signed(25, 9),
    1531 => to_signed(-13, 9),
    1532 => to_signed(-22, 9),
    1533 => to_signed(3, 9),
    1534 => to_signed(2, 9),
    1535 => to_signed(16, 9),
    1536 => to_signed(-11, 9),
    1537 => to_signed(-18, 9),
    1538 => to_signed(10, 9),
    1539 => to_signed(-37, 9),
    1540 => to_signed(-4, 9),
    1541 => to_signed(0, 9),
    1542 => to_signed(2, 9),
    1543 => to_signed(-2, 9),
    1544 => to_signed(-12, 9),
    1545 => to_signed(-18, 9),
    1546 => to_signed(15, 9),
    1547 => to_signed(9, 9),
    1548 => to_signed(-3, 9),
    1549 => to_signed(9, 9),
    1550 => to_signed(42, 9),
    1551 => to_signed(13, 9),
    1552 => to_signed(34, 9),
    1553 => to_signed(68, 9),
    1554 => to_signed(46, 9),
    1555 => to_signed(12, 9),
    1556 => to_signed(2, 9),
    1557 => to_signed(25, 9),
    1558 => to_signed(44, 9),
    1559 => to_signed(37, 9),
    1560 => to_signed(22, 9),
    1561 => to_signed(19, 9),
    1562 => to_signed(0, 9),
    1563 => to_signed(8, 9),
    1564 => to_signed(-1, 9),
    1565 => to_signed(-10, 9),
    1566 => to_signed(-11, 9),
    1567 => to_signed(-28, 9),
    1568 => to_signed(-11, 9),
    1569 => to_signed(-42, 9),
    1570 => to_signed(-23, 9),
    1571 => to_signed(6, 9),
    1572 => to_signed(1, 9),
    1573 => to_signed(-1, 9),
    1574 => to_signed(11, 9),
    1575 => to_signed(3, 9),
    1576 => to_signed(-3, 9),
    1577 => to_signed(-15, 9),
    1578 => to_signed(-12, 9),
    1579 => to_signed(0, 9),
    1580 => to_signed(-3, 9),
    1581 => to_signed(3, 9),
    1582 => to_signed(-17, 9),
    1583 => to_signed(1, 9),
    1584 => to_signed(-21, 9),
    1585 => to_signed(-17, 9),
    1586 => to_signed(3, 9),
    1587 => to_signed(4, 9),
    1588 => to_signed(-2, 9),
    1589 => to_signed(-17, 9),
    1590 => to_signed(-67, 9),
    1591 => to_signed(-42, 9),
    1592 => to_signed(-26, 9),
    1593 => to_signed(-2, 9),
    1594 => to_signed(8, 9),
    1595 => to_signed(0, 9),
    1596 => to_signed(-2, 9),
    1597 => to_signed(-1, 9),
    1598 => to_signed(13, 9),
    1599 => to_signed(-6, 9),
    1600 => to_signed(4, 9),
    1601 => to_signed(0, 9),
    1602 => to_signed(-3, 9),
    1603 => to_signed(-1, 9),
    1604 => to_signed(-2, 9),
    1605 => to_signed(9, 9),
    1606 => to_signed(38, 9),
    1607 => to_signed(35, 9),
    1608 => to_signed(-10, 9),
    1609 => to_signed(-23, 9),
    1610 => to_signed(-13, 9),
    1611 => to_signed(-11, 9),
    1612 => to_signed(7, 9),
    1613 => to_signed(1, 9),
    1614 => to_signed(0, 9),
    1615 => to_signed(-54, 9),
    1616 => to_signed(-23, 9),
    1617 => to_signed(2, 9),
    1618 => to_signed(-2, 9),
    1619 => to_signed(-7, 9),
    1620 => to_signed(-12, 9),
    1621 => to_signed(-16, 9),
    1622 => to_signed(-36, 9),
    1623 => to_signed(-18, 9),
    1624 => to_signed(28, 9),
    1625 => to_signed(3, 9),
    1626 => to_signed(3, 9),
    1627 => to_signed(13, 9),
    1628 => to_signed(17, 9),
    1629 => to_signed(8, 9),
    1630 => to_signed(-4, 9),
    1631 => to_signed(39, 9),
    1632 => to_signed(24, 9),
    1633 => to_signed(4, 9),
    1634 => to_signed(1, 9),
    1635 => to_signed(11, 9),
    1636 => to_signed(14, 9),
    1637 => to_signed(42, 9),
    1638 => to_signed(-5, 9),
    1639 => to_signed(17, 9),
    1640 => to_signed(56, 9),
    1641 => to_signed(-2, 9),
    1642 => to_signed(-3, 9),
    1643 => to_signed(14, 9),
    1644 => to_signed(24, 9),
    1645 => to_signed(-1, 9),
    1646 => to_signed(30, 9),
    1647 => to_signed(33, 9),
    1648 => to_signed(23, 9),
    1649 => to_signed(0, 9),
    1650 => to_signed(3, 9),
    1651 => to_signed(63, 9),
    1652 => to_signed(41, 9),
    1653 => to_signed(14, 9),
    1654 => to_signed(40, 9),
    1655 => to_signed(27, 9),
    1656 => to_signed(-8, 9),
    1657 => to_signed(-2, 9),
    1658 => to_signed(-3, 9),
    1659 => to_signed(49, 9),
    1660 => to_signed(23, 9),
    1661 => to_signed(11, 9),
    1662 => to_signed(-9, 9),
    1663 => to_signed(-10, 9),
    1664 => to_signed(6, 9),
    1665 => to_signed(-2, 9),
    1666 => to_signed(0, 9),
    1667 => to_signed(0, 9),
    1668 => to_signed(-5, 9),
    1669 => to_signed(-34, 9),
    1670 => to_signed(-4, 9),
    1671 => to_signed(-23, 9),
    1672 => to_signed(-9, 9),
    1673 => to_signed(-1, 9),
    1674 => to_signed(2, 9),
    1675 => to_signed(-2, 9),
    1676 => to_signed(2, 9),
    1677 => to_signed(-5, 9),
    1678 => to_signed(1, 9),
    1679 => to_signed(0, 9),
    1680 => to_signed(1, 9),
    1681 => to_signed(3, 9),
    1682 => to_signed(-4, 9),
    1683 => to_signed(-2, 9),
    1684 => to_signed(-1, 9),
    1685 => to_signed(1, 9),
    1686 => to_signed(0, 9),
    1687 => to_signed(-3, 9),
    1688 => to_signed(3, 9),
    1689 => to_signed(-2, 9),
    1690 => to_signed(4, 9),
    1691 => to_signed(-3, 9),
    1692 => to_signed(1, 9),
    1693 => to_signed(1, 9),
    1694 => to_signed(0, 9),
    1695 => to_signed(0, 9),
    1696 => to_signed(-1, 9),
    1697 => to_signed(-1, 9),
    1698 => to_signed(0, 9),
    1699 => to_signed(-4, 9),
    1700 => to_signed(0, 9),
    1701 => to_signed(0, 9),
    1702 => to_signed(-5, 9),
    1703 => to_signed(0, 9),
    1704 => to_signed(-2, 9),
    1705 => to_signed(4, 9),
    1706 => to_signed(-2, 9),
    1707 => to_signed(0, 9),
    1708 => to_signed(-2, 9),
    1709 => to_signed(-2, 9),
    1710 => to_signed(3, 9),
    1711 => to_signed(0, 9),
    1712 => to_signed(0, 9),
    1713 => to_signed(5, 9),
    1714 => to_signed(-1, 9),
    1715 => to_signed(0, 9),
    1716 => to_signed(2, 9),
    1717 => to_signed(-2, 9),
    1718 => to_signed(-2, 9),
    1719 => to_signed(0, 9),
    1720 => to_signed(-3, 9),
    1721 => to_signed(0, 9),
    1722 => to_signed(-2, 9),
    1723 => to_signed(0, 9),
    1724 => to_signed(1, 9),
    1725 => to_signed(2, 9),
    1726 => to_signed(-1, 9),
    1727 => to_signed(-2, 9),
    1728 => to_signed(-5, 9),
    1729 => to_signed(-2, 9),
    1730 => to_signed(-6, 9),
    1731 => to_signed(1, 9),
    1732 => to_signed(-5, 9),
    1733 => to_signed(-4, 9),
    1734 => to_signed(-1, 9),
    1735 => to_signed(0, 9),
    1736 => to_signed(39, 9),
    1737 => to_signed(13, 9),
    1738 => to_signed(-14, 9),
    1739 => to_signed(6, 9),
    1740 => to_signed(12, 9),
    1741 => to_signed(9, 9),
    1742 => to_signed(0, 9),
    1743 => to_signed(4, 9),
    1744 => to_signed(18, 9),
    1745 => to_signed(1, 9),
    1746 => to_signed(-14, 9),
    1747 => to_signed(3, 9),
    1748 => to_signed(5, 9),
    1749 => to_signed(-1, 9),
    1750 => to_signed(0, 9),
    1751 => to_signed(19, 9),
    1752 => to_signed(49, 9),
    1753 => to_signed(22, 9),
    1754 => to_signed(9, 9),
    1755 => to_signed(6, 9),
    1756 => to_signed(-10, 9),
    1757 => to_signed(-2, 9),
    1758 => to_signed(1, 9),
    1759 => to_signed(1, 9),
    1760 => to_signed(21, 9),
    1761 => to_signed(19, 9),
    1762 => to_signed(5, 9),
    1763 => to_signed(26, 9),
    1764 => to_signed(5, 9),
    1765 => to_signed(-2, 9),
    1766 => to_signed(1, 9),
    1767 => to_signed(-9, 9),
    1768 => to_signed(-7, 9),
    1769 => to_signed(-24, 9),
    1770 => to_signed(0, 9),
    1771 => to_signed(-33, 9),
    1772 => to_signed(-18, 9),
    1773 => to_signed(1, 9),
    1774 => to_signed(1, 9),
    1775 => to_signed(11, 9),
    1776 => to_signed(3, 9),
    1777 => to_signed(23, 9),
    1778 => to_signed(11, 9),
    1779 => to_signed(-41, 9),
    1780 => to_signed(-35, 9),
    1781 => to_signed(-4, 9),
    1782 => to_signed(2, 9),
    1783 => to_signed(28, 9),
    1784 => to_signed(12, 9),
    1785 => to_signed(0, 9),
    1786 => to_signed(7, 9),
    1787 => to_signed(-42, 9),
    1788 => to_signed(10, 9),
    1789 => to_signed(4, 9),
    1790 => to_signed(2, 9),
    1791 => to_signed(-5, 9),
    1792 => to_signed(9, 9),
    1793 => to_signed(8, 9),
    1794 => to_signed(-12, 9),
    1795 => to_signed(-11, 9),
    1796 => to_signed(27, 9),
    1797 => to_signed(4, 9),
    1798 => to_signed(26, 9),
    1799 => to_signed(8, 9),
    1800 => to_signed(10, 9),
    1801 => to_signed(41, 9),
    1802 => to_signed(33, 9),
    1803 => to_signed(13, 9),
    1804 => to_signed(3, 9),
    1805 => to_signed(0, 9),
    1806 => to_signed(19, 9),
    1807 => to_signed(51, 9),
    1808 => to_signed(43, 9),
    1809 => to_signed(5, 9),
    1810 => to_signed(-15, 9),
    1811 => to_signed(0, 9),
    1812 => to_signed(-2, 9),
    1813 => to_signed(-11, 9),
    1814 => to_signed(10, 9),
    1815 => to_signed(-1, 9),
    1816 => to_signed(0, 9),
    1817 => to_signed(-24, 9),
    1818 => to_signed(-15, 9),
    1819 => to_signed(0, 9),
    1820 => to_signed(-1, 9),
    1821 => to_signed(4, 9),
    1822 => to_signed(15, 9),
    1823 => to_signed(-25, 9),
    1824 => to_signed(-14, 9),
    1825 => to_signed(21, 9),
    1826 => to_signed(16, 9),
    1827 => to_signed(0, 9),
    1828 => to_signed(2, 9),
    1829 => to_signed(2, 9),
    1830 => to_signed(0, 9),
    1831 => to_signed(-16, 9),
    1832 => to_signed(-11, 9),
    1833 => to_signed(-7, 9),
    1834 => to_signed(19, 9),
    1835 => to_signed(0, 9),
    1836 => to_signed(-5, 9),
    1837 => to_signed(-10, 9),
    1838 => to_signed(-19, 9),
    1839 => to_signed(10, 9),
    1840 => to_signed(-16, 9),
    1841 => to_signed(-21, 9),
    1842 => to_signed(-8, 9),
    1843 => to_signed(-1, 9),
    1844 => to_signed(0, 9),
    1845 => to_signed(-8, 9),
    1846 => to_signed(-6, 9),
    1847 => to_signed(12, 9),
    1848 => to_signed(2, 9),
    1849 => to_signed(-20, 9),
    1850 => to_signed(0, 9),
    1851 => to_signed(4, 9),
    1852 => to_signed(-2, 9),
    1853 => to_signed(0, 9),
    1854 => to_signed(5, 9),
    1855 => to_signed(11, 9),
    1856 => to_signed(-15, 9),
    1857 => to_signed(4, 9),
    1858 => to_signed(11, 9),
    1859 => to_signed(-5, 9),
    1860 => to_signed(-1, 9),
    1861 => to_signed(-2, 9),
    1862 => to_signed(-2, 9),
    1863 => to_signed(0, 9),
    1864 => to_signed(-2, 9),
    1865 => to_signed(0, 9),
    1866 => to_signed(0, 9),
    1867 => to_signed(-4, 9),
    1868 => to_signed(0, 9),
    1869 => to_signed(0, 9),
    1870 => to_signed(0, 9),
    1871 => to_signed(3, 9),
    1872 => to_signed(4, 9),
    1873 => to_signed(0, 9),
    1874 => to_signed(0, 9),
    1875 => to_signed(-2, 9),
    1876 => to_signed(0, 9),
    1877 => to_signed(3, 9),
    1878 => to_signed(1, 9),
    1879 => to_signed(1, 9),
    1880 => to_signed(3, 9),
    1881 => to_signed(-2, 9),
    1882 => to_signed(0, 9),
    1883 => to_signed(-1, 9),
    1884 => to_signed(0, 9),
    1885 => to_signed(-1, 9),
    1886 => to_signed(-3, 9),
    1887 => to_signed(0, 9),
    1888 => to_signed(0, 9),
    1889 => to_signed(-1, 9),
    1890 => to_signed(-4, 9),
    1891 => to_signed(4, 9),
    1892 => to_signed(0, 9),
    1893 => to_signed(2, 9),
    1894 => to_signed(-2, 9),
    1895 => to_signed(0, 9),
    1896 => to_signed(-4, 9),
    1897 => to_signed(1, 9),
    1898 => to_signed(2, 9),
    1899 => to_signed(1, 9),
    1900 => to_signed(-1, 9),
    1901 => to_signed(-4, 9),
    1902 => to_signed(0, 9),
    1903 => to_signed(-1, 9),
    1904 => to_signed(0, 9),
    1905 => to_signed(0, 9),
    1906 => to_signed(-1, 9),
    1907 => to_signed(1, 9),
    1908 => to_signed(0, 9),
    1909 => to_signed(-3, 9),
    1910 => to_signed(1, 9),
    1911 => to_signed(2, 9),
    1912 => to_signed(0, 9),
    1913 => to_signed(-2, 9),
    1914 => to_signed(0, 9),
    1915 => to_signed(-1, 9),
    1916 => to_signed(0, 9),
    1917 => to_signed(-3, 9),
    1918 => to_signed(-3, 9),
    1919 => to_signed(-3, 9),
    1920 => to_signed(6, 9),
    1921 => to_signed(-2, 9),
    1922 => to_signed(7, 9),
    1923 => to_signed(-19, 9),
    1924 => to_signed(19, 9),
    1925 => to_signed(5, 9),
    1926 => to_signed(-2, 9),
    1927 => to_signed(5, 9),
    1928 => to_signed(-5, 9),
    1929 => to_signed(-25, 9),
    1930 => to_signed(-27, 9),
    1931 => to_signed(-1, 9),
    1932 => to_signed(-28, 9),
    1933 => to_signed(-26, 9),
    1934 => to_signed(-14, 9),
    1935 => to_signed(-5, 9),
    1936 => to_signed(4, 9),
    1937 => to_signed(-2, 9),
    1938 => to_signed(19, 9),
    1939 => to_signed(42, 9),
    1940 => to_signed(-6, 9),
    1941 => to_signed(-62, 9),
    1942 => to_signed(-50, 9),
    1943 => to_signed(-2, 9),
    1944 => to_signed(0, 9),
    1945 => to_signed(24, 9),
    1946 => to_signed(41, 9),
    1947 => to_signed(21, 9),
    1948 => to_signed(-28, 9),
    1949 => to_signed(-20, 9),
    1950 => to_signed(12, 9),
    1951 => to_signed(-4, 9),
    1952 => to_signed(-2, 9),
    1953 => to_signed(20, 9),
    1954 => to_signed(15, 9),
    1955 => to_signed(-26, 9),
    1956 => to_signed(-19, 9),
    1957 => to_signed(2, 9),
    1958 => to_signed(39, 9),
    1959 => to_signed(-1, 9),
    1960 => to_signed(0, 9),
    1961 => to_signed(12, 9),
    1962 => to_signed(15, 9),
    1963 => to_signed(24, 9),
    1964 => to_signed(17, 9),
    1965 => to_signed(13, 9),
    1966 => to_signed(30, 9),
    1967 => to_signed(0, 9),
    1968 => to_signed(4, 9),
    1969 => to_signed(7, 9),
    1970 => to_signed(9, 9),
    1971 => to_signed(17, 9),
    1972 => to_signed(22, 9),
    1973 => to_signed(11, 9),
    1974 => to_signed(13, 9),
    1975 => to_signed(0, 9),
    1976 => to_signed(1, 9),
    1977 => to_signed(-5, 9),
    1978 => to_signed(1, 9),
    1979 => to_signed(-10, 9),
    1980 => to_signed(4, 9),
    1981 => to_signed(11, 9),
    1982 => to_signed(2, 9),
    1983 => to_signed(2, 9),
	
    -- biases_L2 (hidden layer biases):
    1984 => to_signed(0, 9),
    1985 => to_signed(0, 9),
    1986 => to_signed(1, 9),
    1987 => to_signed(0, 9),
    1988 => to_signed(0, 9),
    1989 => to_signed(0, 9),
    1990 => to_signed(1, 9),
    1991 => to_signed(-2, 9),
    1992 => to_signed(0, 9),
    1993 => to_signed(0, 9),
    1994 => to_signed(0, 9),
    1995 => to_signed(0, 9),
    1996 => to_signed(0, 9),
    1997 => to_signed(0, 9),
    1998 => to_signed(0, 9),
    1999 => to_signed(0, 9),
    2000 => to_signed(0, 9),
    2001 => to_signed(0, 9),
    2002 => to_signed(0, 9),
    2003 => to_signed(1, 9),
    2004 => to_signed(0, 9),
    2005 => to_signed(0, 9),
    2006 => to_signed(0, 9),
    2007 => to_signed(0, 9),
    2008 => to_signed(-1, 9),
    2009 => to_signed(1, 9),
    2010 => to_signed(2, 9),
    2011 => to_signed(0, 9),
    2012 => to_signed(0, 9),
    2013 => to_signed(0, 9),
    2014 => to_signed(0, 9),
    2015 => to_signed(1, 9),
	
    -- weights_L4 (output layer weights):
    2016 => to_signed(0, 9),
    2017 => to_signed(26, 9),
    2018 => to_signed(-32, 9),
    2019 => to_signed(2, 9),
    2020 => to_signed(26, 9),
    2021 => to_signed(-37, 9),
    2022 => to_signed(107, 9),
    2023 => to_signed(-78, 9),
    2024 => to_signed(-47, 9),
    2025 => to_signed(0, 9),
    2026 => to_signed(2, 9),
    2027 => to_signed(1, 9),
    2028 => to_signed(79, 9),
    2029 => to_signed(-14, 9),
    2030 => to_signed(-32, 9),
    2031 => to_signed(-68, 9),
    2032 => to_signed(0, 9),
    2033 => to_signed(-70, 9),
    2034 => to_signed(-30, 9),
    2035 => to_signed(-21, 9),
    2036 => to_signed(-1, 9),
    2037 => to_signed(-40, 9),
    2038 => to_signed(51, 9),
    2039 => to_signed(-12, 9),
    2040 => to_signed(32, 9),
    2041 => to_signed(-1, 9),
    2042 => to_signed(42, 9),
    2043 => to_signed(1, 9),
    2044 => to_signed(-20, 9),
    2045 => to_signed(18, 9),
    2046 => to_signed(-1, 9),
    2047 => to_signed(10, 9),
    2048 => to_signed(43, 9),
    2049 => to_signed(-109, 9),
    2050 => to_signed(-52, 9),
    2051 => to_signed(-2, 9),
    2052 => to_signed(-18, 9),
    2053 => to_signed(-12, 9),
    2054 => to_signed(-94, 9),
    2055 => to_signed(72, 9),
    2056 => to_signed(21, 9),
    2057 => to_signed(-3, 9),
    2058 => to_signed(3, 9),
    2059 => to_signed(-2, 9),
    2060 => to_signed(4, 9),
    2061 => to_signed(-7, 9),
    2062 => to_signed(55, 9),
    2063 => to_signed(4, 9),
    2064 => to_signed(0, 9),
    2065 => to_signed(58, 9),
    2066 => to_signed(20, 9),
    2067 => to_signed(-41, 9),
    2068 => to_signed(5, 9),
    2069 => to_signed(40, 9),
    2070 => to_signed(-23, 9),
    2071 => to_signed(13, 9),
    2072 => to_signed(94, 9),
    2073 => to_signed(-74, 9),
    2074 => to_signed(-15, 9),
    2075 => to_signed(0, 9),
    2076 => to_signed(21, 9),
    2077 => to_signed(-8, 9),
    2078 => to_signed(2, 9),
    2079 => to_signed(14, 9),
    2080 => to_signed(-56, 9),
    2081 => to_signed(41, 9),
    2082 => to_signed(-78, 9),
    2083 => to_signed(0, 9),
    2084 => to_signed(26, 9),
    2085 => to_signed(23, 9),
    2086 => to_signed(-5, 9),
    2087 => to_signed(58, 9),
    2088 => to_signed(-156, 9),
    2089 => to_signed(-1, 9),
    2090 => to_signed(2, 9),
    2091 => to_signed(26, 9),
    2092 => to_signed(70, 9),
    2093 => to_signed(9, 9),
    2094 => to_signed(28, 9),
    2095 => to_signed(2, 9),
    2096 => to_signed(-6, 9),
    2097 => to_signed(18, 9),
    2098 => to_signed(48, 9),
    2099 => to_signed(-11, 9),
    2100 => to_signed(42, 9),
    2101 => to_signed(20, 9),
    2102 => to_signed(47, 9),
    2103 => to_signed(14, 9),
    2104 => to_signed(-57, 9),
    2105 => to_signed(18, 9),
    2106 => to_signed(-44, 9),
    2107 => to_signed(0, 9),
    2108 => to_signed(31, 9),
    2109 => to_signed(11, 9),
    2110 => to_signed(-2, 9),
    2111 => to_signed(-24, 9),
    2112 => to_signed(-30, 9),
    2113 => to_signed(51, 9),
    2114 => to_signed(-50, 9),
    2115 => to_signed(-2, 9),
    2116 => to_signed(61, 9),
    2117 => to_signed(56, 9),
    2118 => to_signed(-37, 9),
    2119 => to_signed(-4, 9),
    2120 => to_signed(48, 9),
    2121 => to_signed(-4, 9),
    2122 => to_signed(-3, 9),
    2123 => to_signed(13, 9),
    2124 => to_signed(-7, 9),
    2125 => to_signed(65, 9),
    2126 => to_signed(-59, 9),
    2127 => to_signed(77, 9),
    2128 => to_signed(-7, 9),
    2129 => to_signed(24, 9),
    2130 => to_signed(-20, 9),
    2131 => to_signed(7, 9),
    2132 => to_signed(-13, 9),
    2133 => to_signed(24, 9),
    2134 => to_signed(-36, 9),
    2135 => to_signed(0, 9),
    2136 => to_signed(-63, 9),
    2137 => to_signed(44, 9),
    2138 => to_signed(-34, 9),
    2139 => to_signed(0, 9),
    2140 => to_signed(-76, 9),
    2141 => to_signed(-35, 9),
    2142 => to_signed(0, 9),
    2143 => to_signed(-8, 9),
    2144 => to_signed(45, 9),
    2145 => to_signed(-47, 9),
    2146 => to_signed(41, 9),
    2147 => to_signed(-2, 9),
    2148 => to_signed(-107, 9),
    2149 => to_signed(-78, 9),
    2150 => to_signed(20, 9),
    2151 => to_signed(-45, 9),
    2152 => to_signed(13, 9),
    2153 => to_signed(4, 9),
    2154 => to_signed(-4, 9),
    2155 => to_signed(-13, 9),
    2156 => to_signed(-7, 9),
    2157 => to_signed(-24, 9),
    2158 => to_signed(22, 9),
    2159 => to_signed(-58, 9),
    2160 => to_signed(-6, 9),
    2161 => to_signed(48, 9),
    2162 => to_signed(55, 9),
    2163 => to_signed(-3, 9),
    2164 => to_signed(-94, 9),
    2165 => to_signed(37, 9),
    2166 => to_signed(-29, 9),
    2167 => to_signed(-23, 9),
    2168 => to_signed(51, 9),
    2169 => to_signed(-59, 9),
    2170 => to_signed(117, 9),
    2171 => to_signed(-1, 9),
    2172 => to_signed(46, 9),
    2173 => to_signed(-27, 9),
    2174 => to_signed(0, 9),
    2175 => to_signed(80, 9),
    2176 => to_signed(-28, 9),
    2177 => to_signed(-4, 9),
    2178 => to_signed(62, 9),
    2179 => to_signed(0, 9),
    2180 => to_signed(34, 9),
    2181 => to_signed(63, 9),
    2182 => to_signed(32, 9),
    2183 => to_signed(15, 9),
    2184 => to_signed(11, 9),
    2185 => to_signed(1, 9),
    2186 => to_signed(0, 9),
    2187 => to_signed(-3, 9),
    2188 => to_signed(-54, 9),
    2189 => to_signed(-14, 9),
    2190 => to_signed(-34, 9),
    2191 => to_signed(49, 9),
    2192 => to_signed(0, 9),
    2193 => to_signed(-98, 9),
    2194 => to_signed(-24, 9),
    2195 => to_signed(-25, 9),
    2196 => to_signed(-67, 9),
    2197 => to_signed(-81, 9),
    2198 => to_signed(18, 9),
    2199 => to_signed(13, 9),
    2200 => to_signed(10, 9),
    2201 => to_signed(118, 9),
    2202 => to_signed(-95, 9),
    2203 => to_signed(0, 9),
    2204 => to_signed(31, 9),
    2205 => to_signed(66, 9),
    2206 => to_signed(4, 9),
    2207 => to_signed(30, 9),
    2208 => to_signed(65, 9),
    2209 => to_signed(-22, 9),
    2210 => to_signed(12, 9),
    2211 => to_signed(2, 9),
    2212 => to_signed(-19, 9),
    2213 => to_signed(-25, 9),
    2214 => to_signed(9, 9),
    2215 => to_signed(-71, 9),
    2216 => to_signed(-26, 9),
    2217 => to_signed(0, 9),
    2218 => to_signed(1, 9),
    2219 => to_signed(-10, 9),
    2220 => to_signed(-14, 9),
    2221 => to_signed(-4, 9),
    2222 => to_signed(115, 9),
    2223 => to_signed(21, 9),
    2224 => to_signed(13, 9),
    2225 => to_signed(-24, 9),
    2226 => to_signed(66, 9),
    2227 => to_signed(-14, 9),
    2228 => to_signed(18, 9),
    2229 => to_signed(-40, 9),
    2230 => to_signed(56, 9),
    2231 => to_signed(5, 9),
    2232 => to_signed(-40, 9),
    2233 => to_signed(-36, 9),
    2234 => to_signed(-14, 9),
    2235 => to_signed(-1, 9),
    2236 => to_signed(-69, 9),
    2237 => to_signed(-29, 9),
    2238 => to_signed(0, 9),
    2239 => to_signed(40, 9),
    2240 => to_signed(-85, 9),
    2241 => to_signed(-19, 9),
    2242 => to_signed(86, 9),
    2243 => to_signed(1, 9),
    2244 => to_signed(-27, 9),
    2245 => to_signed(18, 9),
    2246 => to_signed(-71, 9),
    2247 => to_signed(-42, 9),
    2248 => to_signed(15, 9),
    2249 => to_signed(0, 9),
    2250 => to_signed(1, 9),
    2251 => to_signed(15, 9),
    2252 => to_signed(-21, 9),
    2253 => to_signed(6, 9),
    2254 => to_signed(0, 9),
    2255 => to_signed(-34, 9),
    2256 => to_signed(1, 9),
    2257 => to_signed(61, 9),
    2258 => to_signed(-36, 9),
    2259 => to_signed(74, 9),
    2260 => to_signed(35, 9),
    2261 => to_signed(108, 9),
    2262 => to_signed(-51, 9),
    2263 => to_signed(-3, 9),
    2264 => to_signed(-52, 9),
    2265 => to_signed(24, 9),
    2266 => to_signed(18, 9),
    2267 => to_signed(-5, 9),
    2268 => to_signed(0, 9),
    2269 => to_signed(55, 9),
    2270 => to_signed(-3, 9),
    2271 => to_signed(-5, 9),
    2272 => to_signed(99, 9),
    2273 => to_signed(10, 9),
    2274 => to_signed(-10, 9),
    2275 => to_signed(-1, 9),
    2276 => to_signed(-3, 9),
    2277 => to_signed(0, 9),
    2278 => to_signed(7, 9),
    2279 => to_signed(48, 9),
    2280 => to_signed(36, 9),
    2281 => to_signed(0, 9),
    2282 => to_signed(-3, 9),
    2283 => to_signed(19, 9),
    2284 => to_signed(-11, 9),
    2285 => to_signed(4, 9),
    2286 => to_signed(-6, 9),
    2287 => to_signed(-3, 9),
    2288 => to_signed(-3, 9),
    2289 => to_signed(-33, 9),
    2290 => to_signed(-21, 9),
    2291 => to_signed(13, 9),
    2292 => to_signed(61, 9),
    2293 => to_signed(-21, 9),
    2294 => to_signed(35, 9),
    2295 => to_signed(-22, 9),
    2296 => to_signed(-15, 9),
    2297 => to_signed(-30, 9),
    2298 => to_signed(19, 9),
    2299 => to_signed(1, 9),
    2300 => to_signed(22, 9),
    2301 => to_signed(-42, 9),
    2302 => to_signed(-3, 9),
    2303 => to_signed(-38, 9),
    2304 => to_signed(-49, 9),
    2305 => to_signed(63, 9),
    2306 => to_signed(34, 9),
    2307 => to_signed(-2, 9),
    2308 => to_signed(14, 9),
    2309 => to_signed(-21, 9),
    2310 => to_signed(37, 9),
    2311 => to_signed(50, 9),
    2312 => to_signed(78, 9),
    2313 => to_signed(2, 9),
    2314 => to_signed(0, 9),
    2315 => to_signed(-38, 9),
    2316 => to_signed(-28, 9),
    2317 => to_signed(-21, 9),
    2318 => to_signed(-79, 9),
    2319 => to_signed(20, 9),
    2320 => to_signed(0, 9),
    2321 => to_signed(24, 9),
    2322 => to_signed(-50, 9),
    2323 => to_signed(18, 9),
    2324 => to_signed(22, 9),
    2325 => to_signed(-48, 9),
    2326 => to_signed(-70, 9),
    2327 => to_signed(3, 9),
    2328 => to_signed(35, 9),
    2329 => to_signed(7, 9),
    2330 => to_signed(0, 9),
    2331 => to_signed(-4, 9),
    2332 => to_signed(13, 9),
    2333 => to_signed(-2, 9),
    2334 => to_signed(0, 9),
    2335 => to_signed(-89, 9),

   -- biases_L4 - 10 adresses (output layer biases):
    2336 => to_signed(-2, 9),
    2337 => to_signed(-8, 9),
    2338 => to_signed(0, 9),
    2339 => to_signed(0, 9),
    2340 => to_signed(8, 9),
    2341 => to_signed(4, 9),
    2342 => to_signed(1, 9),
    2343 => to_signed(1, 9),
    2344 => to_signed(-5, 9),
    2345 => to_signed(1, 9)
);
    
begin
    process(addr)
    begin
        if addr >= 0 and addr <= 2345 then
            data_out <= rom(addr);
        else
            data_out <= (others => '0'); -- Default value for out-of-range address
        end if;
    end process;
end Behavioral;
